* SPICE NETLIST
***************************************

.SUBCKT crtmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT cfmom_mx PLUS1 MINUS1 PLUS2 MINUS2 BULK
.ENDS
***************************************
.SUBCKT lcesd1_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT lcesd2_rf PLUS MINUS
.ENDS
***************************************
.SUBCKT mimcap_2p0_shield PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin TOP BOT
.ENDS
***************************************
.SUBCKT mimcap_2p0_sin_3t PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT mimcap_2p0_wos PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf33_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT moscap_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT nmos_rf D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT nmos_rf33_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmos_rf_6t D G S B NG PG
.ENDS
***************************************
.SUBCKT nmoscap PLUS MINUS
.ENDS
***************************************
.SUBCKT nmoscap_33 PLUS MINUS
.ENDS
***************************************
.SUBCKT pmos_rf D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33 D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf33_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf33_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_5t D G S B PG
.ENDS
***************************************
.SUBCKT pmos_rf_nw D G S B
.ENDS
***************************************
.SUBCKT pmos_rf_nw_5t D G S B PG
.ENDS
***************************************
.SUBCKT rnod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnpo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rnwsti_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpod_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodrpo_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rpodw_m PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1rpo_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppo1w_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_dis PLUS MINUS B
.ENDS
***************************************
.SUBCKT rppolyhri_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolyl_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolys_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT rppolywo_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT sbd_rf_nw PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_std_mu_x_20k PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT spiral_sym_ct_mu_x_20k PLUS MINUS BULK CTAP
.ENDS
***************************************
.SUBCKT spiral_sym_mu_x_20k PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_nr36 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT xjvar_w40 PLUS MINUS BULK
.ENDS
***************************************
.SUBCKT pmos2v_CDNS_6647224192713
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT nmos2v_CDNS_6647224192717
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT MirrorAdder
** N=35 EP=0 IP=18 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: A B Cin VDD GND S Cout
.ENDS
***************************************
.SUBCKT 4bitMirrorAdder GND VDD A2 A3 B0 A0 Cin S0 B1 A1 S1 B2 S2 B3 S3 Cout
** N=67 EP=16 IP=76 FDC=112
M0 27 A0 GND GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=7.695e-13 PD=6.66e-06 PS=3.39e-06 NRD=0.168421 NRS=0.0947368 sa=1.2e-06 sb=4.8e-07 sca=0.435365 scb=1.38069e-08 scc=1.27438e-16 $X=2770 $Y=-18887 $D=0
M1 20 Cin 27 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=1.368e-12 PD=3.39e-06 PS=6.66e-06 NRD=0.0947368 NRS=0.168421 sa=4.8e-07 sb=4.51e-06 sca=0.192279 scb=1.9905e-12 scc=2.1682e-23 $X=5950 $Y=-18887 $D=0
M2 29 B0 20 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=7.695e-13 PD=3.1e-06 PS=3.39e-06 NRD=0.0438596 NRS=0.0947368 sa=1.2e-06 sb=3.79e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=6670 $Y=-18887 $D=0
M3 GND A0 29 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=3.5625e-13 PD=3.39e-06 PS=3.1e-06 NRD=0.0947368 NRS=0.0438596 sa=1.63e-06 sb=3.36e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=7100 $Y=-18887 $D=0
M4 28 B0 GND GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=2.35e-06 sb=2.64e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=7820 $Y=-18887 $D=0
M5 GND A0 28 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=3.07e-06 sb=1.92e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=8540 $Y=-18887 $D=0
M6 28 Cin GND GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=3.79e-06 sb=1.2e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=9260 $Y=-18887 $D=0
M7 30 Cin 21 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=1.368e-12 PD=3.1e-06 PS=6.66e-06 NRD=0.0438596 NRS=0.168421 sa=4.8e-07 sb=1.34e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=12830 $Y=-18887 $D=0
M8 31 B0 30 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=3.5625e-13 PD=3.1e-06 PS=3.1e-06 NRD=0.0438596 NRS=0.0438596 sa=9.1e-07 sb=9.1e-07 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=13260 $Y=-18887 $D=0
M9 GND A0 31 GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=3.5625e-13 PD=6.66e-06 PS=3.1e-06 NRD=0.168421 NRS=0.0438596 sa=1.34e-06 sb=4.8e-07 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=13690 $Y=-18887 $D=0
M10 GND 21 S0 GND N L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.8e-13 PD=1.54e-06 PS=2.96e-06 NRD=0.27 NRS=0.48 sa=4.8e-07 sb=1.2e-06 sca=0.183464 scb=2.64904e-15 scc=1.03277e-29 $X=17360 $Y=-18093 $D=0
M11 3 20 GND GND N L=1.8e-07 W=1e-06 AD=4.8e-13 AS=2.7e-13 PD=2.96e-06 PS=1.54e-06 NRD=0.48 NRS=0.27 sa=1.2e-06 sb=4.8e-07 sca=0.183464 scb=2.64904e-15 scc=1.03277e-29 $X=18080 $Y=-18093 $D=0
M12 GND B0 27 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=1.368e-12 PD=3.39e-06 PS=6.66e-06 NRD=0.0947368 NRS=0.168421 sa=4.8e-07 sb=1.2e-06 sca=0.894508 scb=1.13306e-05 scc=1.39165e-10 $X=2050 $Y=-18887 $D=0
M13 21 20 28 GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=7.695e-13 PD=6.66e-06 PS=3.39e-06 NRD=0.168421 NRS=0.0947368 sa=4.51e-06 sb=4.8e-07 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=9980 $Y=-18887 $D=0
M14 39 A1 GND GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=7.695e-13 PD=6.66e-06 PS=3.39e-06 NRD=0.168421 NRS=0.0947368 sa=1.2e-06 sb=4.8e-07 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=23180 $Y=-18882 $D=0
M15 32 3 39 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=1.368e-12 PD=3.39e-06 PS=6.66e-06 NRD=0.0947368 NRS=0.168421 sa=4.8e-07 sb=4.51e-06 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=26360 $Y=-18882 $D=0
M16 41 B1 32 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=7.695e-13 PD=3.1e-06 PS=3.39e-06 NRD=0.0438596 NRS=0.0947368 sa=1.2e-06 sb=3.79e-06 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=27080 $Y=-18882 $D=0
M17 GND A1 41 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=3.5625e-13 PD=3.39e-06 PS=3.1e-06 NRD=0.0947368 NRS=0.0438596 sa=1.63e-06 sb=3.36e-06 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=27510 $Y=-18882 $D=0
M18 40 B1 GND GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=2.35e-06 sb=2.64e-06 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=28230 $Y=-18882 $D=0
M19 GND A1 40 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=3.07e-06 sb=1.92e-06 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=28950 $Y=-18882 $D=0
M20 40 3 GND GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=3.79e-06 sb=1.2e-06 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=29670 $Y=-18882 $D=0
M21 42 3 33 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=1.368e-12 PD=3.1e-06 PS=6.66e-06 NRD=0.0438596 NRS=0.168421 sa=4.8e-07 sb=1.34e-06 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=33240 $Y=-18882 $D=0
M22 43 B1 42 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=3.5625e-13 PD=3.1e-06 PS=3.1e-06 NRD=0.0438596 NRS=0.0438596 sa=9.1e-07 sb=9.1e-07 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=33670 $Y=-18882 $D=0
M23 GND A1 43 GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=3.5625e-13 PD=6.66e-06 PS=3.1e-06 NRD=0.168421 NRS=0.0438596 sa=1.34e-06 sb=4.8e-07 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=34100 $Y=-18882 $D=0
M24 GND 33 S1 GND N L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.8e-13 PD=1.54e-06 PS=2.96e-06 NRD=0.27 NRS=0.48 sa=4.8e-07 sb=1.2e-06 sca=0.18333 scb=2.52361e-15 scc=9.3591e-30 $X=37770 $Y=-18088 $D=0
M25 4 32 GND GND N L=1.8e-07 W=1e-06 AD=4.8e-13 AS=2.7e-13 PD=2.96e-06 PS=1.54e-06 NRD=0.48 NRS=0.27 sa=1.2e-06 sb=4.8e-07 sca=0.18333 scb=2.52361e-15 scc=9.3591e-30 $X=38490 $Y=-18088 $D=0
M26 GND B1 39 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=1.368e-12 PD=3.39e-06 PS=6.66e-06 NRD=0.0947368 NRS=0.168421 sa=4.8e-07 sb=1.2e-06 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=22460 $Y=-18882 $D=0
M27 33 32 40 GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=7.695e-13 PD=6.66e-06 PS=3.39e-06 NRD=0.168421 NRS=0.0947368 sa=4.51e-06 sb=4.8e-07 sca=0.191745 scb=1.89713e-12 scc=1.96578e-23 $X=30390 $Y=-18882 $D=0
M28 51 A2 GND GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=7.695e-13 PD=6.66e-06 PS=3.39e-06 NRD=0.168421 NRS=0.0947368 sa=1.2e-06 sb=4.8e-07 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=43195 $Y=-18887 $D=0
M29 44 4 51 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=1.368e-12 PD=3.39e-06 PS=6.66e-06 NRD=0.0947368 NRS=0.168421 sa=4.8e-07 sb=4.51e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=46375 $Y=-18887 $D=0
M30 53 B2 44 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=7.695e-13 PD=3.1e-06 PS=3.39e-06 NRD=0.0438596 NRS=0.0947368 sa=1.2e-06 sb=3.79e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=47095 $Y=-18887 $D=0
M31 GND A2 53 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=3.5625e-13 PD=3.39e-06 PS=3.1e-06 NRD=0.0947368 NRS=0.0438596 sa=1.63e-06 sb=3.36e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=47525 $Y=-18887 $D=0
M32 52 B2 GND GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=2.35e-06 sb=2.64e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=48245 $Y=-18887 $D=0
M33 GND A2 52 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=3.07e-06 sb=1.92e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=48965 $Y=-18887 $D=0
M34 52 4 GND GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=3.79e-06 sb=1.2e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=49685 $Y=-18887 $D=0
M35 54 4 45 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=1.368e-12 PD=3.1e-06 PS=6.66e-06 NRD=0.0438596 NRS=0.168421 sa=4.8e-07 sb=1.34e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=53255 $Y=-18887 $D=0
M36 55 B2 54 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=3.5625e-13 PD=3.1e-06 PS=3.1e-06 NRD=0.0438596 NRS=0.0438596 sa=9.1e-07 sb=9.1e-07 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=53685 $Y=-18887 $D=0
M37 GND A2 55 GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=3.5625e-13 PD=6.66e-06 PS=3.1e-06 NRD=0.168421 NRS=0.0438596 sa=1.34e-06 sb=4.8e-07 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=54115 $Y=-18887 $D=0
M38 GND 45 S2 GND N L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.8e-13 PD=1.54e-06 PS=2.96e-06 NRD=0.27 NRS=0.48 sa=4.8e-07 sb=1.2e-06 sca=0.183464 scb=2.64904e-15 scc=1.03277e-29 $X=57785 $Y=-18093 $D=0
M39 6 44 GND GND N L=1.8e-07 W=1e-06 AD=4.8e-13 AS=2.7e-13 PD=2.96e-06 PS=1.54e-06 NRD=0.48 NRS=0.27 sa=1.2e-06 sb=4.8e-07 sca=0.183464 scb=2.64904e-15 scc=1.03277e-29 $X=58505 $Y=-18093 $D=0
M40 GND B2 51 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=1.368e-12 PD=3.39e-06 PS=6.66e-06 NRD=0.0947368 NRS=0.168421 sa=4.8e-07 sb=1.2e-06 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=42475 $Y=-18887 $D=0
M41 45 44 52 GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=7.695e-13 PD=6.66e-06 PS=3.39e-06 NRD=0.168421 NRS=0.0947368 sa=4.51e-06 sb=4.8e-07 sca=0.191897 scb=1.9905e-12 scc=2.1682e-23 $X=50405 $Y=-18887 $D=0
M42 63 A3 GND GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=7.695e-13 PD=6.66e-06 PS=3.39e-06 NRD=0.168421 NRS=0.0947368 sa=1.2e-06 sb=4.8e-07 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=64465 $Y=-18912 $D=0
M43 56 6 63 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=1.368e-12 PD=3.39e-06 PS=6.66e-06 NRD=0.0947368 NRS=0.168421 sa=4.8e-07 sb=4.51e-06 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=67645 $Y=-18912 $D=0
M44 65 B3 56 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=7.695e-13 PD=3.1e-06 PS=3.39e-06 NRD=0.0438596 NRS=0.0947368 sa=1.2e-06 sb=3.79e-06 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=68365 $Y=-18912 $D=0
M45 GND A3 65 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=3.5625e-13 PD=3.39e-06 PS=3.1e-06 NRD=0.0947368 NRS=0.0438596 sa=1.63e-06 sb=3.36e-06 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=68795 $Y=-18912 $D=0
M46 64 B3 GND GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=2.35e-06 sb=2.64e-06 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=69515 $Y=-18912 $D=0
M47 GND A3 64 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=3.07e-06 sb=1.92e-06 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=70235 $Y=-18912 $D=0
M48 64 6 GND GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=7.695e-13 PD=3.39e-06 PS=3.39e-06 NRD=0.0947368 NRS=0.0947368 sa=3.79e-06 sb=1.2e-06 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=70955 $Y=-18912 $D=0
M49 66 6 57 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=1.368e-12 PD=3.1e-06 PS=6.66e-06 NRD=0.0438596 NRS=0.168421 sa=4.8e-07 sb=1.34e-06 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=74525 $Y=-18912 $D=0
M50 67 B3 66 GND N L=1.8e-07 W=2.85e-06 AD=3.5625e-13 AS=3.5625e-13 PD=3.1e-06 PS=3.1e-06 NRD=0.0438596 NRS=0.0438596 sa=9.1e-07 sb=9.1e-07 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=74955 $Y=-18912 $D=0
M51 GND A3 67 GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=3.5625e-13 PD=6.66e-06 PS=3.1e-06 NRD=0.168421 NRS=0.0438596 sa=1.34e-06 sb=4.8e-07 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=75385 $Y=-18912 $D=0
M52 GND 57 S3 GND N L=1.8e-07 W=1e-06 AD=2.7e-13 AS=4.8e-13 PD=1.54e-06 PS=2.96e-06 NRD=0.27 NRS=0.48 sa=4.8e-07 sb=1.2e-06 sca=0.350627 scb=6.28841e-10 scc=2.25438e-19 $X=79055 $Y=-18118 $D=0
M53 Cout 56 GND GND N L=1.8e-07 W=1e-06 AD=4.8e-13 AS=2.7e-13 PD=2.96e-06 PS=1.54e-06 NRD=0.48 NRS=0.27 sa=1.2e-06 sb=4.8e-07 sca=0.59762 scb=5.64653e-07 scc=2.69942e-13 $X=79775 $Y=-18118 $D=0
M54 GND B3 63 GND N L=1.8e-07 W=2.85e-06 AD=7.695e-13 AS=1.368e-12 PD=3.39e-06 PS=6.66e-06 NRD=0.0947368 NRS=0.168421 sa=4.8e-07 sb=1.2e-06 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=63745 $Y=-18912 $D=0
M55 57 56 64 GND N L=1.8e-07 W=2.85e-06 AD=1.368e-12 AS=7.695e-13 PD=6.66e-06 PS=3.39e-06 NRD=0.168421 NRS=0.0947368 sa=4.51e-06 sb=4.8e-07 sca=0.192678 scb=2.53083e-12 scc=3.53905e-23 $X=71675 $Y=-18912 $D=0
M56 22 A0 VDD VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=1.215e-12 PD=9.96e-06 PS=5.04e-06 NRD=0.106667 NRS=0.06 sa=1.2e-06 sb=4.8e-07 sca=0.776587 scb=8.26593e-05 scc=2.31282e-07 $X=2770 $Y=-11615 $D=16
M57 20 Cin 22 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=2.16e-12 PD=5.04e-06 PS=9.96e-06 NRD=0.06 NRS=0.106667 sa=4.8e-07 sb=4.51e-06 sca=0.532073 scb=8.26448e-05 scc=2.31282e-07 $X=5950 $Y=-11615 $D=16
M58 23 B0 20 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=1.215e-12 PD=4.75e-06 PS=5.04e-06 NRD=0.0277778 NRS=0.06 sa=1.2e-06 sb=3.79e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=6670 $Y=-11615 $D=16
M59 VDD A0 23 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=5.625e-13 PD=5.04e-06 PS=4.75e-06 NRD=0.06 NRS=0.0277778 sa=1.63e-06 sb=3.36e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=7100 $Y=-11615 $D=16
M60 24 B0 VDD VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=2.35e-06 sb=2.64e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=7820 $Y=-11615 $D=16
M61 VDD A0 24 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=3.07e-06 sb=1.92e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=8540 $Y=-11615 $D=16
M62 24 Cin VDD VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=3.79e-06 sb=1.2e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=9260 $Y=-11615 $D=16
M63 25 Cin 21 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=2.16e-12 PD=4.75e-06 PS=9.96e-06 NRD=0.0277778 NRS=0.106667 sa=4.8e-07 sb=1.34e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=12830 $Y=-11615 $D=16
M64 26 A0 25 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=5.625e-13 PD=4.75e-06 PS=4.75e-06 NRD=0.0277778 NRS=0.0277778 sa=9.1e-07 sb=9.1e-07 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=13260 $Y=-11615 $D=16
M65 VDD B0 26 VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=5.625e-13 PD=9.96e-06 PS=4.75e-06 NRD=0.106667 NRS=0.0277778 sa=1.34e-06 sb=4.8e-07 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=13690 $Y=-11615 $D=16
M66 VDD 21 S0 VDD P L=1.8e-07 W=1.5e-06 AD=4.05e-13 AS=7.2e-13 PD=2.04e-06 PS=3.96e-06 NRD=0.18 NRS=0.32 sa=4.8e-07 sb=1.2e-06 sca=0.927846 scb=0.000131515 scc=1.75553e-07 $X=17360 $Y=-11540 $D=16
M67 3 20 VDD VDD P L=1.8e-07 W=1.5e-06 AD=7.2e-13 AS=4.05e-13 PD=3.96e-06 PS=2.04e-06 NRD=0.32 NRS=0.18 sa=1.2e-06 sb=4.8e-07 sca=0.927846 scb=0.000131515 scc=1.75553e-07 $X=18080 $Y=-11540 $D=16
M68 VDD B0 22 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=2.16e-12 PD=5.04e-06 PS=9.96e-06 NRD=0.06 NRS=0.106667 sa=4.8e-07 sb=1.2e-06 sca=1.24067 scb=9.4504e-05 scc=2.31435e-07 $X=2050 $Y=-11615 $D=16
M69 21 20 24 VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=1.215e-12 PD=9.96e-06 PS=5.04e-06 NRD=0.106667 NRS=0.06 sa=4.51e-06 sb=4.8e-07 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=9980 $Y=-11615 $D=16
M70 34 A1 VDD VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=1.215e-12 PD=9.96e-06 PS=5.04e-06 NRD=0.106667 NRS=0.06 sa=1.2e-06 sb=4.8e-07 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=23180 $Y=-11610 $D=16
M71 32 3 34 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=2.16e-12 PD=5.04e-06 PS=9.96e-06 NRD=0.06 NRS=0.106667 sa=4.8e-07 sb=4.51e-06 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=26360 $Y=-11610 $D=16
M72 35 B1 32 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=1.215e-12 PD=4.75e-06 PS=5.04e-06 NRD=0.0277778 NRS=0.06 sa=1.2e-06 sb=3.79e-06 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=27080 $Y=-11610 $D=16
M73 VDD A1 35 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=5.625e-13 PD=5.04e-06 PS=4.75e-06 NRD=0.06 NRS=0.0277778 sa=1.63e-06 sb=3.36e-06 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=27510 $Y=-11610 $D=16
M74 36 B1 VDD VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=2.35e-06 sb=2.64e-06 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=28230 $Y=-11610 $D=16
M75 VDD A1 36 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=3.07e-06 sb=1.92e-06 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=28950 $Y=-11610 $D=16
M76 36 3 VDD VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=3.79e-06 sb=1.2e-06 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=29670 $Y=-11610 $D=16
M77 37 3 33 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=2.16e-12 PD=4.75e-06 PS=9.96e-06 NRD=0.0277778 NRS=0.106667 sa=4.8e-07 sb=1.34e-06 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=33240 $Y=-11610 $D=16
M78 38 A1 37 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=5.625e-13 PD=4.75e-06 PS=4.75e-06 NRD=0.0277778 NRS=0.0277778 sa=9.1e-07 sb=9.1e-07 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=33670 $Y=-11610 $D=16
M79 VDD B1 38 VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=5.625e-13 PD=9.96e-06 PS=4.75e-06 NRD=0.106667 NRS=0.0277778 sa=1.34e-06 sb=4.8e-07 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=34100 $Y=-11610 $D=16
M80 VDD 33 S1 VDD P L=1.8e-07 W=1.5e-06 AD=4.05e-13 AS=7.2e-13 PD=2.04e-06 PS=3.96e-06 NRD=0.18 NRS=0.32 sa=4.8e-07 sb=1.2e-06 sca=0.918954 scb=0.000126014 scc=1.60097e-07 $X=37770 $Y=-11535 $D=16
M81 4 32 VDD VDD P L=1.8e-07 W=1.5e-06 AD=7.2e-13 AS=4.05e-13 PD=3.96e-06 PS=2.04e-06 NRD=0.32 NRS=0.18 sa=1.2e-06 sb=4.8e-07 sca=0.918954 scb=0.000126014 scc=1.60097e-07 $X=38490 $Y=-11535 $D=16
M82 VDD B1 34 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=2.16e-12 PD=5.04e-06 PS=9.96e-06 NRD=0.06 NRS=0.106667 sa=4.8e-07 sb=1.2e-06 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=22460 $Y=-11610 $D=16
M83 33 32 36 VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=1.215e-12 PD=9.96e-06 PS=5.04e-06 NRD=0.106667 NRS=0.06 sa=4.51e-06 sb=4.8e-07 sca=0.52761 scb=7.92585e-05 scc=2.11141e-07 $X=30390 $Y=-11610 $D=16
M84 46 A2 VDD VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=1.215e-12 PD=9.96e-06 PS=5.04e-06 NRD=0.106667 NRS=0.06 sa=1.2e-06 sb=4.8e-07 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=43195 $Y=-11615 $D=16
M85 44 4 46 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=2.16e-12 PD=5.04e-06 PS=9.96e-06 NRD=0.06 NRS=0.106667 sa=4.8e-07 sb=4.51e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=46375 $Y=-11615 $D=16
M86 47 B2 44 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=1.215e-12 PD=4.75e-06 PS=5.04e-06 NRD=0.0277778 NRS=0.06 sa=1.2e-06 sb=3.79e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=47095 $Y=-11615 $D=16
M87 VDD A2 47 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=5.625e-13 PD=5.04e-06 PS=4.75e-06 NRD=0.06 NRS=0.0277778 sa=1.63e-06 sb=3.36e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=47525 $Y=-11615 $D=16
M88 48 B2 VDD VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=2.35e-06 sb=2.64e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=48245 $Y=-11615 $D=16
M89 VDD A2 48 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=3.07e-06 sb=1.92e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=48965 $Y=-11615 $D=16
M90 48 4 VDD VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=3.79e-06 sb=1.2e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=49685 $Y=-11615 $D=16
M91 49 4 45 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=2.16e-12 PD=4.75e-06 PS=9.96e-06 NRD=0.0277778 NRS=0.106667 sa=4.8e-07 sb=1.34e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=53255 $Y=-11615 $D=16
M92 50 A2 49 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=5.625e-13 PD=4.75e-06 PS=4.75e-06 NRD=0.0277778 NRS=0.0277778 sa=9.1e-07 sb=9.1e-07 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=53685 $Y=-11615 $D=16
M93 VDD B2 50 VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=5.625e-13 PD=9.96e-06 PS=4.75e-06 NRD=0.106667 NRS=0.0277778 sa=1.34e-06 sb=4.8e-07 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=54115 $Y=-11615 $D=16
M94 VDD 45 S2 VDD P L=1.8e-07 W=1.5e-06 AD=4.05e-13 AS=7.2e-13 PD=2.04e-06 PS=3.96e-06 NRD=0.18 NRS=0.32 sa=4.8e-07 sb=1.2e-06 sca=0.927846 scb=0.000131515 scc=1.75553e-07 $X=57785 $Y=-11540 $D=16
M95 6 44 VDD VDD P L=1.8e-07 W=1.5e-06 AD=7.2e-13 AS=4.05e-13 PD=3.96e-06 PS=2.04e-06 NRD=0.32 NRS=0.18 sa=1.2e-06 sb=4.8e-07 sca=0.927846 scb=0.000131515 scc=1.75553e-07 $X=58505 $Y=-11540 $D=16
M96 VDD B2 46 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=2.16e-12 PD=5.04e-06 PS=9.96e-06 NRD=0.06 NRS=0.106667 sa=4.8e-07 sb=1.2e-06 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=42475 $Y=-11615 $D=16
M97 45 44 48 VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=1.215e-12 PD=9.96e-06 PS=5.04e-06 NRD=0.106667 NRS=0.06 sa=4.51e-06 sb=4.8e-07 sca=0.531614 scb=8.26448e-05 scc=2.31282e-07 $X=50405 $Y=-11615 $D=16
M98 58 A3 VDD VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=1.215e-12 PD=9.96e-06 PS=5.04e-06 NRD=0.106667 NRS=0.06 sa=1.2e-06 sb=4.8e-07 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=64465 $Y=-11640 $D=16
M99 56 6 58 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=2.16e-12 PD=5.04e-06 PS=9.96e-06 NRD=0.06 NRS=0.106667 sa=4.8e-07 sb=4.51e-06 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=67645 $Y=-11640 $D=16
M100 59 B3 56 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=1.215e-12 PD=4.75e-06 PS=5.04e-06 NRD=0.0277778 NRS=0.06 sa=1.2e-06 sb=3.79e-06 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=68365 $Y=-11640 $D=16
M101 VDD A3 59 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=5.625e-13 PD=5.04e-06 PS=4.75e-06 NRD=0.06 NRS=0.0277778 sa=1.63e-06 sb=3.36e-06 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=68795 $Y=-11640 $D=16
M102 60 B3 VDD VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=2.35e-06 sb=2.64e-06 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=69515 $Y=-11640 $D=16
M103 VDD A3 60 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=3.07e-06 sb=1.92e-06 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=70235 $Y=-11640 $D=16
M104 60 6 VDD VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=1.215e-12 PD=5.04e-06 PS=5.04e-06 NRD=0.06 NRS=0.06 sa=3.79e-06 sb=1.2e-06 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=70955 $Y=-11640 $D=16
M105 61 6 57 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=2.16e-12 PD=4.75e-06 PS=9.96e-06 NRD=0.0277778 NRS=0.106667 sa=4.8e-07 sb=1.34e-06 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=74525 $Y=-11640 $D=16
M106 62 A3 61 VDD P L=1.8e-07 W=4.5e-06 AD=5.625e-13 AS=5.625e-13 PD=4.75e-06 PS=4.75e-06 NRD=0.0277778 NRS=0.0277778 sa=9.1e-07 sb=9.1e-07 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=74955 $Y=-11640 $D=16
M107 VDD B3 62 VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=5.625e-13 PD=9.96e-06 PS=4.75e-06 NRD=0.106667 NRS=0.0277778 sa=1.34e-06 sb=4.8e-07 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=75385 $Y=-11640 $D=16
M108 VDD 57 S3 VDD P L=1.8e-07 W=1.5e-06 AD=4.05e-13 AS=7.2e-13 PD=2.04e-06 PS=3.96e-06 NRD=0.18 NRS=0.32 sa=4.8e-07 sb=1.2e-06 sca=1.21681 scb=0.000162719 scc=2.78042e-07 $X=79055 $Y=-11565 $D=16
M109 Cout 56 VDD VDD P L=1.8e-07 W=1.5e-06 AD=7.2e-13 AS=4.05e-13 PD=3.96e-06 PS=2.04e-06 NRD=0.32 NRS=0.18 sa=1.2e-06 sb=4.8e-07 sca=1.67109 scb=0.000173531 scc=2.78168e-07 $X=79775 $Y=-11565 $D=16
M110 VDD B3 58 VDD P L=1.8e-07 W=4.5e-06 AD=1.215e-12 AS=2.16e-12 PD=5.04e-06 PS=9.96e-06 NRD=0.06 NRS=0.106667 sa=4.8e-07 sb=1.2e-06 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=63745 $Y=-11640 $D=16
M111 57 56 60 VDD P L=1.8e-07 W=4.5e-06 AD=2.16e-12 AS=1.215e-12 PD=9.96e-06 PS=5.04e-06 NRD=0.106667 NRS=0.06 sa=4.51e-06 sb=4.8e-07 sca=0.552953 scb=0.000101769 scc=3.64296e-07 $X=71675 $Y=-11640 $D=16
.ENDS
***************************************
